** Profile: "SCHEMATIC1-Vout"  [ D:\altele\Etti\OrcadCIS lite proiecte\SERS_Petre_Adrian\SERS_Petre_Adrian_432E-PSpiceFiles\SCHEMATIC1\Vout.sim ] 

** Creating circuit file "Vout.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "d:/altele/etti/spice models/draghici/lib_modelepspice_anexa_1/modele_a1_lib/bzx84c2v7.lib" 
.LIB "d:/altele/aplicatii/cadence/tools/capture/library/pspice/modele_a1_lib/mjd31cg.lib" 
.LIB "d:/altele/aplicatii/cadence/tools/capture/library/pspice/modele_a1_lib/bc846b.lib" 
.LIB "d:/altele/aplicatii/cadence/tools/capture/library/pspice/modele_a1_lib/bzx84c5v1.lib" 
.LIB "d:/altele/aplicatii/cadence/tools/capture/library/pspice/modele_a1_lib/bc856b.lib" 
* From [PSPICE NETLIST] section of C:\Users\adria\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V1 0 50 5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
